// tb.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module tb (
	);

	wire         resize_inst_resized_image_valid;                                                          // resize_inst:resized_image_valid -> stream_sink_dpi_bfm_resize_resized_image_inst:sink_valid
	wire  [31:0] resize_inst_resized_image_data;                                                           // resize_inst:resized_image_data -> stream_sink_dpi_bfm_resize_resized_image_inst:sink_data
	wire         resize_inst_resized_image_ready;                                                          // stream_sink_dpi_bfm_resize_resized_image_inst:sink_ready -> resize_inst:resized_image_ready
	wire         stream_source_dpi_bfm_resize_original_image_inst_source_valid;                            // stream_source_dpi_bfm_resize_original_image_inst:source_valid -> resize_inst:original_image_valid
	wire  [31:0] stream_source_dpi_bfm_resize_original_image_inst_source_data;                             // stream_source_dpi_bfm_resize_original_image_inst:source_data -> resize_inst:original_image_data
	wire         stream_source_dpi_bfm_resize_original_image_inst_source_ready;                            // resize_inst:original_image_ready -> stream_source_dpi_bfm_resize_original_image_inst:source_ready
	wire         clock_reset_inst_clock_clk;                                                               // clock_reset_inst:clock -> [component_dpi_controller_resize_inst:clock, irq_mapper:clk, main_dpi_controller_inst:clock, resize_inst:clock, stream_sink_dpi_bfm_resize_resized_image_inst:clock, stream_source_dpi_bfm_resize_cols_inst:clock, stream_source_dpi_bfm_resize_original_image_inst:clock, stream_source_dpi_bfm_resize_ratio_inst:clock, stream_source_dpi_bfm_resize_rows_inst:clock]
	wire         clock_reset_inst_clock2x_clk;                                                             // clock_reset_inst:clock2x -> [component_dpi_controller_resize_inst:clock2x, main_dpi_controller_inst:clock2x, stream_sink_dpi_bfm_resize_resized_image_inst:clock2x, stream_source_dpi_bfm_resize_cols_inst:clock2x, stream_source_dpi_bfm_resize_original_image_inst:clock2x, stream_source_dpi_bfm_resize_ratio_inst:clock2x, stream_source_dpi_bfm_resize_rows_inst:clock2x]
	wire         component_dpi_controller_resize_inst_component_call_valid;                                // component_dpi_controller_resize_inst:start -> resize_inst:start
	wire         resize_inst_call_stall;                                                                   // resize_inst:busy -> component_dpi_controller_resize_inst:busy
	wire         component_dpi_controller_resize_inst_component_done_conduit;                              // component_dpi_controller_resize_inst:component_done -> concatenate_component_done_inst:in_conduit_0
	wire   [0:0] main_dpi_controller_inst_component_enabled_conduit;                                       // main_dpi_controller_inst:component_enabled -> split_component_start_inst:in_conduit
	wire         component_dpi_controller_resize_inst_component_wait_for_stream_writes_conduit;            // component_dpi_controller_resize_inst:component_wait_for_stream_writes -> concatenate_component_wait_for_stream_writes_inst:in_conduit_0
	wire         component_dpi_controller_resize_inst_dpi_control_bind_conduit;                            // component_dpi_controller_resize_inst:bind_interfaces -> resize_component_dpi_controller_bind_conduit_fanout_inst:in_conduit
	wire         component_dpi_controller_resize_inst_dpi_control_enable_conduit;                          // component_dpi_controller_resize_inst:enable_interfaces -> resize_component_dpi_controller_enable_conduit_fanout_inst:in_conduit
	wire         stream_sink_dpi_bfm_resize_resized_image_inst_dpi_control_stream_active_conduit;          // stream_sink_dpi_bfm_resize_resized_image_inst:stream_active -> resize_component_dpi_controller_stream_active_concatenate_inst:in_conduit_0
	wire         concatenate_component_done_inst_out_conduit_conduit;                                      // concatenate_component_done_inst:out_conduit -> main_dpi_controller_inst:component_done
	wire         concatenate_component_wait_for_stream_writes_inst_out_conduit_conduit;                    // concatenate_component_wait_for_stream_writes_inst:out_conduit -> main_dpi_controller_inst:component_wait_for_stream_writes
	wire         resize_component_dpi_controller_stream_active_concatenate_inst_out_conduit_conduit;       // resize_component_dpi_controller_stream_active_concatenate_inst:out_conduit -> component_dpi_controller_resize_inst:stream_writes_active
	wire         split_component_start_inst_out_conduit_0_conduit;                                         // split_component_start_inst:out_conduit_0 -> component_dpi_controller_resize_inst:component_enabled
	wire         resize_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit;           // resize_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_0 -> stream_source_dpi_bfm_resize_cols_inst:do_bind
	wire         resize_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit;         // resize_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_0 -> stream_source_dpi_bfm_resize_cols_inst:enable
	wire         resize_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit; // resize_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_0 -> stream_source_dpi_bfm_resize_cols_inst:source_ready
	wire         resize_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit;           // resize_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_1 -> stream_source_dpi_bfm_resize_original_image_inst:do_bind
	wire         resize_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit;         // resize_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_1 -> stream_source_dpi_bfm_resize_original_image_inst:enable
	wire         resize_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit; // resize_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_1 -> stream_source_dpi_bfm_resize_ratio_inst:source_ready
	wire         resize_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_2_conduit;           // resize_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_2 -> stream_source_dpi_bfm_resize_ratio_inst:do_bind
	wire         resize_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_2_conduit;         // resize_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_2 -> stream_source_dpi_bfm_resize_ratio_inst:enable
	wire         resize_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_2_conduit; // resize_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_2 -> stream_source_dpi_bfm_resize_rows_inst:source_ready
	wire         resize_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_3_conduit;           // resize_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_3 -> stream_sink_dpi_bfm_resize_resized_image_inst:do_bind
	wire         resize_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_3_conduit;         // resize_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_3 -> stream_sink_dpi_bfm_resize_resized_image_inst:enable
	wire         resize_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_4_conduit;           // resize_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_4 -> stream_source_dpi_bfm_resize_rows_inst:do_bind
	wire         resize_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_4_conduit;         // resize_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_4 -> stream_source_dpi_bfm_resize_rows_inst:enable
	wire         component_dpi_controller_resize_inst_read_implicit_streams_conduit;                       // component_dpi_controller_resize_inst:read_implicit_streams -> resize_component_dpi_controller_implicit_ready_conduit_fanout_inst:in_conduit
	wire         main_dpi_controller_inst_reset_ctrl_conduit;                                              // main_dpi_controller_inst:trigger_reset -> clock_reset_inst:trigger_reset
	wire         resize_inst_return_valid;                                                                 // resize_inst:done -> component_dpi_controller_resize_inst:done
	wire         component_dpi_controller_resize_inst_component_return_stall;                              // component_dpi_controller_resize_inst:stall -> resize_inst:stall
	wire  [31:0] stream_source_dpi_bfm_resize_cols_inst_source_data_data;                                  // stream_source_dpi_bfm_resize_cols_inst:source_data -> resize_inst:cols
	wire  [31:0] stream_source_dpi_bfm_resize_ratio_inst_source_data_data;                                 // stream_source_dpi_bfm_resize_ratio_inst:source_data -> resize_inst:ratio
	wire  [31:0] stream_source_dpi_bfm_resize_rows_inst_source_data_data;                                  // stream_source_dpi_bfm_resize_rows_inst:source_data -> resize_inst:rows
	wire         clock_reset_inst_reset_reset;                                                             // clock_reset_inst:resetn -> [component_dpi_controller_resize_inst:resetn, irq_mapper:reset, main_dpi_controller_inst:resetn, resize_inst:resetn, stream_sink_dpi_bfm_resize_resized_image_inst:resetn, stream_source_dpi_bfm_resize_cols_inst:resetn, stream_source_dpi_bfm_resize_original_image_inst:resetn, stream_source_dpi_bfm_resize_ratio_inst:resetn, stream_source_dpi_bfm_resize_rows_inst:resetn]
	wire         component_dpi_controller_resize_inst_component_irq_irq;                                   // irq_mapper:sender_irq -> component_dpi_controller_resize_inst:done_irq

	hls_sim_clock_reset #(
		.RESET_CYCLE_HOLD (4)
	) clock_reset_inst (
		.clock         (clock_reset_inst_clock_clk),                  //      clock.clk
		.resetn        (clock_reset_inst_reset_reset),                //      reset.reset_n
		.clock2x       (clock_reset_inst_clock2x_clk),                //    clock2x.clk
		.trigger_reset (main_dpi_controller_inst_reset_ctrl_conduit)  // reset_ctrl.conduit
	);

	hls_sim_component_dpi_controller #(
		.COMPONENT_NAME               ("resize"),
		.RETURN_DATAWIDTH             (64),
		.COMPONENT_NUM_SLAVES         (0),
		.COMPONENT_HAS_SLAVE_RETURN   (0),
		.COMPONENT_NUM_OUTPUT_STREAMS (1)
	) component_dpi_controller_resize_inst (
		.clock                            (clock_reset_inst_clock_clk),                                                         //                            clock.clk
		.resetn                           (clock_reset_inst_reset_reset),                                                       //                            reset.reset_n
		.clock2x                          (clock_reset_inst_clock2x_clk),                                                       //                          clock2x.clk
		.bind_interfaces                  (component_dpi_controller_resize_inst_dpi_control_bind_conduit),                      //                 dpi_control_bind.conduit
		.enable_interfaces                (component_dpi_controller_resize_inst_dpi_control_enable_conduit),                    //               dpi_control_enable.conduit
		.stream_writes_active             (resize_component_dpi_controller_stream_active_concatenate_inst_out_conduit_conduit), // dpi_control_stream_writes_active.conduit
		.component_enabled                (split_component_start_inst_out_conduit_0_conduit),                                   //                component_enabled.conduit
		.component_done                   (component_dpi_controller_resize_inst_component_done_conduit),                        //                   component_done.conduit
		.component_wait_for_stream_writes (component_dpi_controller_resize_inst_component_wait_for_stream_writes_conduit),      // component_wait_for_stream_writes.conduit
		.read_implicit_streams            (component_dpi_controller_resize_inst_read_implicit_streams_conduit),                 //            read_implicit_streams.conduit
		.readback_from_slaves             (),                                                                                   //             readback_from_slaves.conduit
		.start                            (component_dpi_controller_resize_inst_component_call_valid),                          //                   component_call.valid
		.busy                             (resize_inst_call_stall),                                                             //                                 .stall
		.done                             (resize_inst_return_valid),                                                           //                 component_return.valid
		.stall                            (component_dpi_controller_resize_inst_component_return_stall),                        //                                 .stall
		.done_irq                         (component_dpi_controller_resize_inst_component_irq_irq),                             //                    component_irq.irq
		.returndata                       ()                                                                                    //                       returndata.data
	);

	tb_concatenate_component_done_inst concatenate_component_done_inst (
		.out_conduit  (concatenate_component_done_inst_out_conduit_conduit),         //  out_conduit.conduit
		.in_conduit_0 (component_dpi_controller_resize_inst_component_done_conduit)  // in_conduit_0.conduit
	);

	tb_concatenate_component_done_inst concatenate_component_wait_for_stream_writes_inst (
		.out_conduit  (concatenate_component_wait_for_stream_writes_inst_out_conduit_conduit),         //  out_conduit.conduit
		.in_conduit_0 (component_dpi_controller_resize_inst_component_wait_for_stream_writes_conduit)  // in_conduit_0.conduit
	);

	hls_sim_main_dpi_controller #(
		.NUM_COMPONENTS                    (1),
		.COMPONENT_NAMES_STR               ("resize"),
		.SIM_COMPONENT_CALL_COUNT_LOG_FILE (".")
	) main_dpi_controller_inst (
		.clock                            (clock_reset_inst_clock_clk),                                            //                            clock.clk
		.resetn                           (clock_reset_inst_reset_reset),                                          //                            reset.reset_n
		.clock2x                          (clock_reset_inst_clock2x_clk),                                          //                          clock2x.clk
		.component_enabled                (main_dpi_controller_inst_component_enabled_conduit),                    //                component_enabled.conduit
		.component_done                   (concatenate_component_done_inst_out_conduit_conduit),                   //                   component_done.conduit
		.component_wait_for_stream_writes (concatenate_component_wait_for_stream_writes_inst_out_conduit_conduit), // component_wait_for_stream_writes.conduit
		.trigger_reset                    (main_dpi_controller_inst_reset_ctrl_conduit)                            //                       reset_ctrl.conduit
	);

	tb_resize_component_dpi_controller_bind_conduit_fanout_inst resize_component_dpi_controller_bind_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_resize_inst_dpi_control_bind_conduit),                  //    in_conduit.conduit
		.out_conduit_0 (resize_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit), // out_conduit_0.conduit
		.out_conduit_1 (resize_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit), // out_conduit_1.conduit
		.out_conduit_2 (resize_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_2_conduit), // out_conduit_2.conduit
		.out_conduit_3 (resize_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_3_conduit), // out_conduit_3.conduit
		.out_conduit_4 (resize_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_4_conduit)  // out_conduit_4.conduit
	);

	tb_resize_component_dpi_controller_bind_conduit_fanout_inst resize_component_dpi_controller_enable_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_resize_inst_dpi_control_enable_conduit),                  //    in_conduit.conduit
		.out_conduit_0 (resize_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit), // out_conduit_0.conduit
		.out_conduit_1 (resize_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit), // out_conduit_1.conduit
		.out_conduit_2 (resize_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_2_conduit), // out_conduit_2.conduit
		.out_conduit_3 (resize_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_3_conduit), // out_conduit_3.conduit
		.out_conduit_4 (resize_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_4_conduit)  // out_conduit_4.conduit
	);

	tb_resize_component_dpi_controller_implicit_ready_conduit_fanout_inst resize_component_dpi_controller_implicit_ready_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_resize_inst_read_implicit_streams_conduit),                       //    in_conduit.conduit
		.out_conduit_0 (resize_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit), // out_conduit_0.conduit
		.out_conduit_1 (resize_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit), // out_conduit_1.conduit
		.out_conduit_2 (resize_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_2_conduit)  // out_conduit_2.conduit
	);

	tb_concatenate_component_done_inst resize_component_dpi_controller_stream_active_concatenate_inst (
		.out_conduit  (resize_component_dpi_controller_stream_active_concatenate_inst_out_conduit_conduit), //  out_conduit.conduit
		.in_conduit_0 (stream_sink_dpi_bfm_resize_resized_image_inst_dpi_control_stream_active_conduit)     // in_conduit_0.conduit
	);

	tb_resize_inst resize_inst (
		.start                (component_dpi_controller_resize_inst_component_call_valid),     //           call.valid
		.busy                 (resize_inst_call_stall),                                        //               .stall
		.clock                (clock_reset_inst_clock_clk),                                    //          clock.clk
		.cols                 (stream_source_dpi_bfm_resize_cols_inst_source_data_data),       //           cols.data
		.original_image_data  (stream_source_dpi_bfm_resize_original_image_inst_source_data),  // original_image.data
		.original_image_ready (stream_source_dpi_bfm_resize_original_image_inst_source_ready), //               .ready
		.original_image_valid (stream_source_dpi_bfm_resize_original_image_inst_source_valid), //               .valid
		.ratio                (stream_source_dpi_bfm_resize_ratio_inst_source_data_data),      //          ratio.data
		.resetn               (clock_reset_inst_reset_reset),                                  //          reset.reset_n
		.resized_image_data   (resize_inst_resized_image_data),                                //  resized_image.data
		.resized_image_ready  (resize_inst_resized_image_ready),                               //               .ready
		.resized_image_valid  (resize_inst_resized_image_valid),                               //               .valid
		.done                 (resize_inst_return_valid),                                      //         return.valid
		.stall                (component_dpi_controller_resize_inst_component_return_stall),   //               .stall
		.rows                 (stream_source_dpi_bfm_resize_rows_inst_source_data_data)        //           rows.data
	);

	tb_split_component_start_inst split_component_start_inst (
		.in_conduit    (main_dpi_controller_inst_component_enabled_conduit), //    in_conduit.conduit
		.out_conduit_0 (split_component_start_inst_out_conduit_0_conduit)    // out_conduit_0.conduit
	);

	hls_sim_stream_sink_dpi_bfm #(
		.COMPONENT_NAME   ("resize"),
		.INTERFACE_NAME   ("resized_image"),
		.STREAM_DATAWIDTH (32),
		.READY_LATENCY    (0)
	) stream_sink_dpi_bfm_resize_resized_image_inst (
		.clock              (clock_reset_inst_clock_clk),                                                       //                     clock.clk
		.resetn             (clock_reset_inst_reset_reset),                                                     //                     reset.reset_n
		.clock2x            (clock_reset_inst_clock2x_clk),                                                     //                   clock2x.clk
		.do_bind            (resize_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_3_conduit),   //          dpi_control_bind.conduit
		.enable             (resize_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_3_conduit), //        dpi_control_enable.conduit
		.stream_active      (stream_sink_dpi_bfm_resize_resized_image_inst_dpi_control_stream_active_conduit),  // dpi_control_stream_active.conduit
		.sink_data          (resize_inst_resized_image_data),                                                   //                      sink.data
		.sink_ready         (resize_inst_resized_image_ready),                                                  //                          .ready
		.sink_valid         (resize_inst_resized_image_valid),                                                  //                          .valid
		.sink_startofpacket (1'b0),                                                                             //               (terminated)
		.sink_endofpacket   (1'b0)                                                                              //               (terminated)
	);

	hls_sim_stream_source_dpi_bfm #(
		.COMPONENT_NAME   ("resize"),
		.INTERFACE_NAME   ("cols"),
		.STREAM_DATAWIDTH (32)
	) stream_source_dpi_bfm_resize_cols_inst (
		.clock        (clock_reset_inst_clock_clk),                                                               //              clock.clk
		.resetn       (clock_reset_inst_reset_reset),                                                             //              reset.reset_n
		.clock2x      (clock_reset_inst_clock2x_clk),                                                             //            clock2x.clk
		.do_bind      (resize_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit),           //   dpi_control_bind.conduit
		.enable       (resize_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit),         // dpi_control_enable.conduit
		.source_data  (stream_source_dpi_bfm_resize_cols_inst_source_data_data),                                  //        source_data.data
		.source_ready (resize_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit), //       source_ready.conduit
		.source_valid ()                                                                                          //             source.conduit
	);

	hls_sim_stream_source_dpi_bfm #(
		.COMPONENT_NAME   ("resize"),
		.INTERFACE_NAME   ("original_image"),
		.STREAM_DATAWIDTH (32)
	) stream_source_dpi_bfm_resize_original_image_inst (
		.clock        (clock_reset_inst_clock_clk),                                                       //              clock.clk
		.resetn       (clock_reset_inst_reset_reset),                                                     //              reset.reset_n
		.clock2x      (clock_reset_inst_clock2x_clk),                                                     //            clock2x.clk
		.do_bind      (resize_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit),   //   dpi_control_bind.conduit
		.enable       (resize_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit), // dpi_control_enable.conduit
		.source_data  (stream_source_dpi_bfm_resize_original_image_inst_source_data),                     //             source.data
		.source_ready (stream_source_dpi_bfm_resize_original_image_inst_source_ready),                    //                   .ready
		.source_valid (stream_source_dpi_bfm_resize_original_image_inst_source_valid)                     //                   .valid
	);

	hls_sim_stream_source_dpi_bfm #(
		.COMPONENT_NAME   ("resize"),
		.INTERFACE_NAME   ("ratio"),
		.STREAM_DATAWIDTH (32)
	) stream_source_dpi_bfm_resize_ratio_inst (
		.clock        (clock_reset_inst_clock_clk),                                                               //              clock.clk
		.resetn       (clock_reset_inst_reset_reset),                                                             //              reset.reset_n
		.clock2x      (clock_reset_inst_clock2x_clk),                                                             //            clock2x.clk
		.do_bind      (resize_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_2_conduit),           //   dpi_control_bind.conduit
		.enable       (resize_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_2_conduit),         // dpi_control_enable.conduit
		.source_data  (stream_source_dpi_bfm_resize_ratio_inst_source_data_data),                                 //        source_data.data
		.source_ready (resize_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit), //       source_ready.conduit
		.source_valid ()                                                                                          //             source.conduit
	);

	hls_sim_stream_source_dpi_bfm #(
		.COMPONENT_NAME   ("resize"),
		.INTERFACE_NAME   ("rows"),
		.STREAM_DATAWIDTH (32)
	) stream_source_dpi_bfm_resize_rows_inst (
		.clock        (clock_reset_inst_clock_clk),                                                               //              clock.clk
		.resetn       (clock_reset_inst_reset_reset),                                                             //              reset.reset_n
		.clock2x      (clock_reset_inst_clock2x_clk),                                                             //            clock2x.clk
		.do_bind      (resize_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_4_conduit),           //   dpi_control_bind.conduit
		.enable       (resize_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_4_conduit),         // dpi_control_enable.conduit
		.source_data  (stream_source_dpi_bfm_resize_rows_inst_source_data_data),                                  //        source_data.data
		.source_ready (resize_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_2_conduit), //       source_ready.conduit
		.source_valid ()                                                                                          //             source.conduit
	);

	tb_irq_mapper irq_mapper (
		.clk        (clock_reset_inst_clock_clk),                             //       clk.clk
		.reset      (~clock_reset_inst_reset_reset),                          // clk_reset.reset
		.sender_irq (component_dpi_controller_resize_inst_component_irq_irq)  //    sender.irq
	);

endmodule
